module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 ;
  assign n61 = ( x9 & x10 ) | ( x9 & x11 ) | ( x10 & x11 ) ;
  assign n62 = x10 ^ x9 ^ 1'b0 ;
  assign n63 = ( x11 & n61 ) | ( x11 & n62 ) | ( n61 & n62 ) ;
  assign n64 = ( ~x12 & x13 ) | ( ~x12 & n63 ) | ( x13 & n63 ) ;
  assign n65 = n64 ^ x12 ^ 1'b0 ;
  assign n66 = ( x12 & n64 ) | ( x12 & n65 ) | ( n64 & n65 ) ;
  assign n67 = n66 ^ x14 ^ 1'b0 ;
  assign n68 = x14 & n66 ;
  assign n69 = x15 & n68 ;
  assign n70 = x16 | n69 ;
  assign n71 = n70 ^ x17 ^ 1'b0 ;
  assign n72 = x17 & n70 ;
  assign n73 = x18 | n72 ;
  assign n74 = x19 & n73 ;
  assign n75 = x20 & n74 ;
  assign n76 = x21 | n75 ;
  assign n77 = n76 ^ x22 ^ 1'b0 ;
  assign n78 = x22 | n76 ;
  assign n79 = x23 & n78 ;
  assign n80 = x24 & n79 ;
  assign n81 = x25 & n80 ;
  assign n82 = x26 | n81 ;
  assign n83 = n82 ^ x27 ^ 1'b0 ;
  assign n84 = x27 & n82 ;
  assign n85 = n84 ^ x28 ^ 1'b0 ;
  assign n86 = ( x9 & x29 ) | ( x9 & n85 ) | ( x29 & n85 ) ;
  assign n87 = ~x9 & n86 ;
  assign n88 = n83 & n87 ;
  assign n89 = n80 ^ x25 ^ 1'b0 ;
  assign n90 = ( x26 & n88 ) | ( x26 & n89 ) | ( n88 & n89 ) ;
  assign n91 = ~x26 & n90 ;
  assign n92 = n78 ^ x23 ^ 1'b0 ;
  assign n93 = n79 ^ x24 ^ 1'b0 ;
  assign n94 = n92 & n93 ;
  assign n95 = n91 & n94 ;
  assign n96 = ~n77 & n95 ;
  assign n97 = n74 ^ x20 ^ 1'b0 ;
  assign n98 = ( x21 & n96 ) | ( x21 & n97 ) | ( n96 & n97 ) ;
  assign n99 = ~x21 & n98 ;
  assign n100 = n72 ^ x18 ^ 1'b0 ;
  assign n101 = n73 ^ x19 ^ 1'b0 ;
  assign n102 = ~n100 & n101 ;
  assign n103 = n99 & n102 ;
  assign n104 = n71 & n103 ;
  assign n105 = n68 ^ x15 ^ 1'b0 ;
  assign n106 = ( x16 & n104 ) | ( x16 & n105 ) | ( n104 & n105 ) ;
  assign n107 = ~x16 & n106 ;
  assign n108 = n67 & n107 ;
  assign n109 = ~n65 & n108 ;
  assign n110 = n61 ^ x11 ^ 1'b0 ;
  assign n111 = n109 & n110 ;
  assign n112 = x7 & x8 ;
  assign n113 = n111 & n112 ;
  assign n114 = x5 & x6 ;
  assign n115 = n113 & n114 ;
  assign n116 = x3 & x4 ;
  assign n117 = n115 & n116 ;
  assign n118 = x1 & x2 ;
  assign n119 = n117 & n118 ;
  assign n120 = x0 & n119 ;
  assign n121 = x28 & x29 ;
  assign n122 = n84 & n121 ;
  assign n123 = n120 | n122 ;
  assign n124 = x1 | x2 ;
  assign n125 = x3 | x4 ;
  assign n126 = n124 | n125 ;
  assign n127 = x5 | x6 ;
  assign n128 = n126 | n127 ;
  assign n129 = x7 | x8 ;
  assign n130 = n128 | n129 ;
  assign n131 = ( x11 & n62 ) | ( x11 & n130 ) | ( n62 & n130 ) ;
  assign n132 = ~n130 & n131 ;
  assign n133 = n63 ^ x12 ^ 1'b0 ;
  assign n134 = ( x13 & n132 ) | ( x13 & n133 ) | ( n132 & n133 ) ;
  assign n135 = ~x13 & n134 ;
  assign n136 = ~n67 & n135 ;
  assign n137 = ( ~x15 & x16 ) | ( ~x15 & n68 ) | ( x16 & n68 ) ;
  assign n138 = n137 ^ n68 ^ 1'b0 ;
  assign n139 = n136 & n138 ;
  assign n140 = ~n71 & n100 ;
  assign n141 = n139 & n140 ;
  assign n142 = ~n101 & n141 ;
  assign n143 = ( ~x20 & x21 ) | ( ~x20 & n74 ) | ( x21 & n74 ) ;
  assign n144 = n143 ^ n74 ^ 1'b0 ;
  assign n145 = n142 & n144 ;
  assign n146 = n77 & n145 ;
  assign n147 = ~n92 & n146 ;
  assign n148 = ~n93 & n147 ;
  assign n149 = ( ~x25 & x26 ) | ( ~x25 & n80 ) | ( x26 & n80 ) ;
  assign n150 = n149 ^ n80 ^ 1'b0 ;
  assign n151 = n148 & n150 ;
  assign n152 = ~n83 & n151 ;
  assign n153 = ~n85 & n152 ;
  assign n154 = x9 & n153 ;
  assign n155 = n122 & ~n154 ;
  assign n156 = n123 & ~n155 ;
  assign n157 = ( x39 & x40 ) | ( x39 & x41 ) | ( x40 & x41 ) ;
  assign n158 = x40 ^ x39 ^ 1'b0 ;
  assign n159 = ( x41 & n157 ) | ( x41 & n158 ) | ( n157 & n158 ) ;
  assign n160 = ( ~x42 & x43 ) | ( ~x42 & n159 ) | ( x43 & n159 ) ;
  assign n161 = n160 ^ x42 ^ 1'b0 ;
  assign n162 = ( x42 & n160 ) | ( x42 & n161 ) | ( n160 & n161 ) ;
  assign n163 = x44 & n162 ;
  assign n164 = x45 & n163 ;
  assign n165 = x46 | n164 ;
  assign n166 = x47 & n165 ;
  assign n167 = x48 | n166 ;
  assign n168 = x49 & n167 ;
  assign n169 = x50 & n168 ;
  assign n170 = x51 | n169 ;
  assign n171 = x52 | n170 ;
  assign n172 = x53 & n171 ;
  assign n173 = x54 & n172 ;
  assign n174 = x55 & n173 ;
  assign n175 = x56 | n174 ;
  assign n176 = x57 & n175 ;
  assign n177 = x58 & x59 ;
  assign n178 = n176 & n177 ;
  assign n179 = x0 & ~n178 ;
  assign n180 = n162 ^ x44 ^ 1'b0 ;
  assign n181 = n165 ^ x47 ^ 1'b0 ;
  assign n182 = n170 ^ x52 ^ 1'b0 ;
  assign n183 = n175 ^ x57 ^ 1'b0 ;
  assign n184 = n176 ^ x58 ^ 1'b0 ;
  assign n185 = x30 & ~x39 ;
  assign n186 = x59 & n185 ;
  assign n187 = n184 & n186 ;
  assign n188 = n183 & n187 ;
  assign n189 = n173 ^ x55 ^ 1'b0 ;
  assign n190 = ( x56 & n188 ) | ( x56 & n189 ) | ( n188 & n189 ) ;
  assign n191 = ~x56 & n190 ;
  assign n192 = n171 ^ x53 ^ 1'b0 ;
  assign n193 = n172 ^ x54 ^ 1'b0 ;
  assign n194 = n192 & n193 ;
  assign n195 = n191 & n194 ;
  assign n196 = ~n182 & n195 ;
  assign n197 = n168 ^ x50 ^ 1'b0 ;
  assign n198 = ( x51 & n196 ) | ( x51 & n197 ) | ( n196 & n197 ) ;
  assign n199 = ~x51 & n198 ;
  assign n200 = n166 ^ x48 ^ 1'b0 ;
  assign n201 = n167 ^ x49 ^ 1'b0 ;
  assign n202 = ~n200 & n201 ;
  assign n203 = n199 & n202 ;
  assign n204 = n181 & n203 ;
  assign n205 = n163 ^ x45 ^ 1'b0 ;
  assign n206 = ( x46 & n204 ) | ( x46 & n205 ) | ( n204 & n205 ) ;
  assign n207 = ~x46 & n206 ;
  assign n208 = n180 & n207 ;
  assign n209 = ~n161 & n208 ;
  assign n210 = n157 ^ x41 ^ 1'b0 ;
  assign n211 = n209 & n210 ;
  assign n212 = x37 & x38 ;
  assign n213 = n211 & n212 ;
  assign n214 = x35 & x36 ;
  assign n215 = n213 & n214 ;
  assign n216 = x33 & x34 ;
  assign n217 = n215 & n216 ;
  assign n218 = x31 & x32 ;
  assign n219 = n217 & n218 ;
  assign n220 = x0 | x30 ;
  assign n221 = x31 | x32 ;
  assign n222 = x33 | x34 ;
  assign n223 = n221 | n222 ;
  assign n224 = x35 | x36 ;
  assign n225 = n223 | n224 ;
  assign n226 = x37 | x38 ;
  assign n227 = n225 | n226 ;
  assign n228 = ( x41 & n158 ) | ( x41 & n227 ) | ( n158 & n227 ) ;
  assign n229 = ~n227 & n228 ;
  assign n230 = n159 ^ x42 ^ 1'b0 ;
  assign n231 = ( x43 & n229 ) | ( x43 & n230 ) | ( n229 & n230 ) ;
  assign n232 = ~x43 & n231 ;
  assign n233 = ~n180 & n232 ;
  assign n234 = ( ~x45 & x46 ) | ( ~x45 & n163 ) | ( x46 & n163 ) ;
  assign n235 = n234 ^ n163 ^ 1'b0 ;
  assign n236 = n233 & n235 ;
  assign n237 = ~n181 & n200 ;
  assign n238 = n236 & n237 ;
  assign n239 = ~n201 & n238 ;
  assign n240 = ( ~x50 & x51 ) | ( ~x50 & n168 ) | ( x51 & n168 ) ;
  assign n241 = n240 ^ n168 ^ 1'b0 ;
  assign n242 = n239 & n241 ;
  assign n243 = n182 & n242 ;
  assign n244 = ~n192 & n243 ;
  assign n245 = ~n193 & n244 ;
  assign n246 = ( ~x55 & x56 ) | ( ~x55 & n173 ) | ( x56 & n173 ) ;
  assign n247 = n246 ^ n173 ^ 1'b0 ;
  assign n248 = n245 & n247 ;
  assign n249 = ~n183 & n248 ;
  assign n250 = ~n184 & n249 ;
  assign n251 = x39 & n250 ;
  assign n252 = ~n220 & n251 ;
  assign n253 = n178 | n252 ;
  assign n254 = ( n219 & ~n252 ) | ( n219 & n253 ) | ( ~n252 & n253 ) ;
  assign n255 = n123 & n254 ;
  assign n256 = ~n179 & n255 ;
  assign n257 = n155 | n256 ;
  assign n258 = x0 & x30 ;
  assign n259 = n251 | n258 ;
  assign n260 = ( n178 & n258 ) | ( n178 & ~n259 ) | ( n258 & ~n259 ) ;
  assign n261 = n156 & n260 ;
  assign y0 = ~n156 ;
  assign y1 = ~n257 ;
  assign y2 = n261 ;
  assign y3 = 1'b0 ;
  assign y4 = 1'b0 ;
  assign y5 = 1'b0 ;
  assign y6 = 1'b0 ;
  assign y7 = 1'b0 ;
  assign y8 = 1'b0 ;
  assign y9 = 1'b0 ;
  assign y10 = 1'b0 ;
  assign y11 = 1'b0 ;
  assign y12 = 1'b0 ;
  assign y13 = 1'b0 ;
  assign y14 = 1'b0 ;
  assign y15 = 1'b0 ;
  assign y16 = 1'b0 ;
  assign y17 = 1'b0 ;
  assign y18 = 1'b0 ;
  assign y19 = 1'b0 ;
  assign y20 = 1'b0 ;
  assign y21 = 1'b0 ;
  assign y22 = 1'b0 ;
  assign y23 = 1'b0 ;
  assign y24 = 1'b0 ;
  assign y25 = 1'b0 ;
  assign y26 = 1'b0 ;
  assign y27 = 1'b0 ;
  assign y28 = 1'b0 ;
  assign y29 = 1'b0 ;
endmodule
